`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:20:28 06/08/2021 
// Design Name: 
// Module Name:    AlU_Control 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module AlU_Control(
    input [1:0] Alu_op ,
    input [5:0] F_Field,
    output [3:0] Operation
    );


endmodule
